module hazard_detection(

//input previous instruction pipeline regwrite flag
//input previous instruction pipeline destination register
//input ex/mem alu data lines


);

endmodule 